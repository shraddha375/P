module matrix_add(a, b, c);
 input [15:0] a;
 input [15:0] b;
 output [15:0] c;

 assign c = a + b; 
 
endmodule
